module PE(

// Input
input Clock
input rst_n

// Input controll signal
input data_clear
input en_shift_right
input en_shift_bottom

input [15:0] b_reg
input b_we

// Output
output [15:0] a_shift_to_righit
output [15:0] partial_sum_to_bottom

TBD
) {

TBD

}
